module Vr8inprior3(I, A, IDLE);
  input [7:0] I;
  output reg [2:0] A;
  output reg IDLE;

  /* Your code below */
endmodule