module Vr7seg (DIG, EN, SEGA, SEGB, SEGC, SEGD, SEGE, SEGF, SEGG);
  input [3:0] DIG;
  input EN;
  output reg SEGA, SEGB, SEGC, SEGD, SEGE, SEGF, SEGG;
  reg [1:7] SEGS;

  /* Your code below */ 
endmodule
